module test_control();

endmodule